PK   G�~S�8��  �.    cirkitFile.json��oɕ�����*u���d /��"/�� �fF�F�R�L����[���[-�}�36�� ���>�xX��CV��e�_�4�������i�?���-�Zq��a����~���j���?��ۯ?��x���yy��a�����>_��ͪL��mYn��m��몼^vî�t�z��]���x�����+XX!�f�*��3DR_��
���Q���a��B�0CT!��0CT!�m�!���.�U�5*^(��(��Zi�b���r����������������������s�x�Kd�x�Kd
`���E�v�%2E�v�%2E�v�%2E�v�%2E�v�%2E�v�%2E�v�%r&��ΰD���ΰD���ΰD� bz�v������������������������H}��a�L��a�L��a�L��a�L|���U�v�%2E�v�%2E�v�%2E�v�%2E�v�%R_�kgX"S�kgX"Sx��,����a�ܯon/O#������������E���p]>{F��?~�����-Wi�[��jWo���Y�u��EgE��]�	�Kx/�a�LQFS|����?���AX"S�?��"�q��񏃰D���AX"S�?��">�I�-)��Y� ��*&g,������Z�|2�vcmG錥K}�zW�ޡt�ҥ�d�+Y�Ft_���C�Oc�Xc��k;Jg,]����լw(��ty��zװޡt�ҥ~�z�b�C錥K}�zײޡt�ҥ�c��X�P:c�|y%<����g0�/����	�L�hbp618��|��b\�?8��|��2b�?8i�|��h�?8m�|���m�?8q�|���s�?8u�|��ry�?8y�|��B�?8}�|����i8�|���
�?8�|����?����8p�(������[q`���1�{��n����t�r�l�հ�-7U7,S���v�ViU�)���|�l=]X>{��_J��_����S�g0�o���S�g0_z�.�N=,�x�ӷ�W-����M,��|�7^��&��`>�U	��&��`>�
��&��`>��
�G�*�C��{pa������织a���������a�������;�a�������{�a��������a���������Y�*8�|�yg�?8�|�yO�?8�|�y7�?8�|�y�?z{
�?��?*8�|�y��?8�|�y��?8�|�y��?8�|�y��?8�|�y�ֿ�,��|����,��|�(��?X>�����?X>���	��?X>���}��E��#��5�?X>������?X>���A��?X>������?X>���)�_���`>o'����`�4�^I�!���>�}U�Og��f��:o�8���.�3/?o_8������{�ź���� I���Y���7]�y�y�ԙ����.�"�軺�<��H���߇�c��^|'����{�y�����蠷�ן���{�yg޹u88�F�ͽ>8�F��ͽ>8�Fwͽ>8�F�eͽ>8�FT�� ��ѡP��_Y[\�nٔ͐�w�,�bU-��F������Y�E�}z�_t��ؿpk�P���ǅ�0�(�%3�'������Ǉ��կ�o���������,��^�(��Y�$t<y�!����3D���Tv�:���AB��"H�x~;C	Osg� ����$t:�*�\���6V�+ܔ��Lx�	�݆oJ�t^<Ą�o�
8�t:Kb�j�aE�R:�31au���8�t:�b������V�)��i�V���SJ���!&��X��N��CLX/�:N)��w�P��x��qJ)�����oR��R�:^bu�R��V�K��SJ�ac��x��qJ�;`LX��:N)��u�	��V�)%�Y�1q߉s_�cu���8��j1&��WX��|�'Ƅ��
�㔒�R�~���x��qJ�؞�����LX�O��RjVA&���X���k}�ҟ�0au���8��;~0&���X��|g
Ƅ���㔒����:�`��)��;%�7����	��IXGk�_����������m7�
V����|#�
��`5	k:�?«���Y��*��y� \�U�j�<��z�V�q@�j�<G��z�n�q@�j�ԟ7 �UA_�&aM�yc\�U�j�ԟ7,�UA_�&a�5��`�I\Z����f����%�]��e��e��%�5��5�x�I_Z����y���&�5����x�IaZ������$&�5����x�IcZ�������D&�5���x�IeZ�����\&�5��U�x��eZ����+���_�D?�irY��e�&�IhMC�F=c���cZ�'G	mz���V��$��N@к�B��
M.�К���Vj���2	�ih}���[M.���˴@M��B��$����=���I�\&�5��=�x��eZ���j���\&�5���x+Z���eZ�Ӯ�V��$������o5�LBkZ�1��V��$����^	o5�LBkZ����V��$�����o5�LBkZ��!���2	�ih����[M.�К��{�h���2	�ih����[M.�К��{�h��$m%��J��*M.�К��{i���2	�ih����[M.�К��{8i���2	�ih���[M.�К��{jI��5�LBkZ���V��$����go5�LBkZ�զ�V��$�����so5�LBkZ�V��C��C��jM.�5�LBkZ�e��V��$������o5�LBkZ�-��V��$�����oM.�К��{}j���2	�ih�g��[M.{��اs���':��T��M;��vDe���L�����W��T��=Se���L��~ԳO�*]v��c@���yԵ}/3z�}�+Ìߩ�U��Lt{�+��3G��L�A�+3ѹ|n�cF����se�Q<uJ�\fO�9W��S'.ΕaF�Թ�s?u�Q<uz�g����uQ�M�y��6˶XU�v�m���]9|yVs�
���7�E*_|?u��Uզ[��f����n���a�R���m�V�ɗ��#�ؗ�F�Of�e��}�pX���_>��?������xدo���?� JG�"H(�G� �t�$�� !���1O D�P:f�Jǜ�AB阙"H(�B	�S�cJ$W�����m�
7��N��a�j�aśRJ�0�0a�۰N)�S�g��nX�����	��V�)�t�j�a������V�)�t��a��x��qJ)���b��:^`u�RJ�o�&��X�����<&�cu���8��p0&�����X���c	Ƅ���㔒w����:^bu�R�V�+��SJ� c��x��qJ�w�cL�w�ܗ�X��:N)��`�	��V�)%߉�1au���8��;��~�:^cu�R�vV�k��SJ��c�~��~���x��qJ�w�`LX��:N)���	��V�)%�a�1au����������(��iQ?�jV���~��V}U���5��](�*諂�$��u�UA_�&a͹K��)  �$�y$�u� q@�j�<G��:j�8�`5	k�G� hU�W�IXS?�@���*XM�Q Z�U�jV_�	��%�5��m�x+J]�إ�]�	^�I^Z���Zs����%�5����x�I`Z�������&�5��a�x�IbZ���^���4&�5��)�x�IdZ�������T&�5��������eZ���^%���\&�5���x+�EL���&��\Vhr���4��N�&�IhMC�{�4�jr���4��'Q�&�IhMC�{+5�jr���4��GT�&�IhMC�{]5�jr���4��gW�0I��$������o5�LBkZ�C��V��$������oE�E�5����R��$������o5�LBkZ�1��V��$����^	o5�LBkZ����V��$�����o5�LBkZ��!���2	�ih����[M.�К��{�h���2	�ih����[M.�К��{�h��$m%��J��*M.�К��{i���2	�ih����[M.�К��{8i���2	�ih���[M.�К��{jI��5�LBkZ���V��$����go5�LBkZ�զ�V��$�����so5�LBkZ�V��C��C��jM.�5�LBkZ�e��V��$������o5�LBkZ�-��V��$�����oM.�К��{}j���2	�ih�g��[M.���e�3O��t;Se�7������>�3U&:o�T��=Se���L��~�3U&:H�T���<w�A���S��Εa���Ѫse�<u��\fO:W��S�qΕ�j03��N��+Ì⩳ ��0�x��Ź2�(�:�p�.3��N�,����.�ݲ)�!ϕ�f��j��mW�C�+�/�j.RaX����H��n����t�r�l�հ�-7U7,S�а�Ҫ��/�|ї�T����U�������}����ms���f?<�n��ö������a�x��]`V������W_ORc$���|�):��G߭���L�_φ{�x��
=�:�s6�Co��y3�F.R�2��Jo���o�v�c��@��\(^���|��%4�[�DPR�����?͚�Ï�?�i��n���]��wF��=Ԅӓ����~�	����ے�8f�)�EC�~���7~}/x��z�����׼�RN�χ����3����닯8��T¯��3���Y�Ԥ������ۅ�o���AOٲ!yi�~��d�8�=|�����8����o���N���Ǜ���/�A����qeq�t�(H�H�ߑ�a�t�}.H�H�UKA��D:�z
R�%�q�T�",�����a�t\��K�㪯 EX"�V�E�Q=��	�O
h\#��E9�j@�k��һ(PG(�q�tZ�� j��4��N��@=-�z�H��Qb>JLH�zZ �4��Nk8�@=-�z�H�U�Q��@=�k��:�(PO���5�i%m4J���i\�{�D�'">POK���5��7�����q�#p ���i\��@=��z�� PO+���5��*�A|gJ|i
��
��q�i	p ���i\�{%@=��z��|���@=��z�8�@�v���S���Z�c�"�T���q�㚴�=e(�5P|���	� �o߸�78��� �7��Mi ��6�dv�1��̨Q�w���-�#�N|g�4��&���DA;GM��O��3�/���C���g0_:_hL�!�����}��v,n�.���>�A;Y>�����o��5�|Y>���,�oԯ5�|Y>��R?j���!��|�~�~��C�c��K���*�������K��4�O`B�	}�&�!J�TB��s���&4�З����&4�З��҉&4�З'�ҩ&4�ЗV���&4�З����&4�З���	&4�З���)&4�з��[�9&4�зA��9&4�зp��?�࿠�9��sJA���h�4�1�
2��~�Zq���tl9�L���-c³ר	:@���N10�ф����N10�ф�Y��C:����NC�/D�
�PSС&4����ыI�PM�{i�PM��(i�PM�{@i�at��	}�*�!j`B�	}�-�!�b`B�	}�0�![`B�	}�3�![`B�	}�6�![`B�	}�9�!�S`B�	}�<�aE���hB��O{H���hB�O@{H���hB�@{H���hB�A{�o[����9��sJE���hB��A{H���hB�%B{H���hB�B{H���hB��B{H���hB�?{X�9&4��{���9&4������9&4�Л��9&4��;*��9&4�лA��[��=�tN��R�9&4���n��9&4��[���9&4��۝��9&4��[��6tN�	�&�6s��tN�	�&L���QA���k�9c�/ �<Js�=q�����3�u+�y������v_��7�H�׻�͔�>�y��g��VGO��uc�"2�7:z�'�������lsF}~�
D�������sF�l�V��H�5W :Ǉc�����qTs�#q| �\��H�4��0:Ǉ}XY[\�nٔ͐g(m�l�U�lw۶+�ݕ�k3����>�+o����}p�Iܯo�}���;g��'��W��27[?�;�?��ޗ����w�4�L�?�}��[�|���������s��������5������n~�̯(����W~E�W~E�W~E�W~E�W�q�>?���?_X]�zו��n�'�E����.�i5\o6ih��:_��y���"_��n7E���m��V�a�n�b���UovE�\>�2���n8��џt4e}����N�Cy�,%��,W���~�����`��|xT>��ϫг�_ �����<c���udĵ��:�i&`.�����Y~L��Ѕ���-<�v����v�n�荫��?����ǵ�x��o*>�T�o*?�T�o�>�T�o�?�T�oj>�ԌoZ}�i基����ɘ������7Q.2�)�������/��}�"���v����m=��������������f8N*~�p���a��x8�o�ܭ�?��W��ַ���?Í|���ċ�_?����wʺ�����Ðo|��y������~��Ǜ��]�=d�l����������<�������� �(y��n��e[�Y�WE]����N��|�<��n�*��U]��J��I�f�n��7�zUU>��L���x�%����&�F����C��������U{��R���S]�]�s���-��k��k��k��klꚢ���h&o�'�ʳkV��RS���k������s�t����[��klꚲ���l'�i&��'�)'�)��y��tK;z}>�2~M?�2~M?�2~M?�2~M?�2~M?���k근?���~s������������N�7�Mʕ?Z�������n�xs��_~���WG��7Gg���	_\5e}�j˓��Ӣ�ˑn��^�(5��f�Y��v���6m���n8/������T?�l쮚�#���</�[}�ּ|�湚�^�����O�:�i���Vm�X�uWEY��κ�nʶ�U�<}!�vX���^��`��Z/�mιEW�:O9�M�:!.J�_~!�g�ݛT�ڪ��}�To�i���;�|�lkR}��,��*ϗw�ݲ��z����]U}�l/������6W����ҳ��y�j�F������KwC�P����j���\5WE���٠:��es���蛕�z���PK   ؚ~Sk2��XP  �Q  /   images/0deaa9e5-55e1-404a-9dfe-2921a303d637.png̛�s%���'�I&�mMl�N&�ļ�Ķm�Ƙ؞$۶m��}���MW���u��?{���p%I8\�o߾!HK��|���u���vA��~���*-&��[��&o1������)�8E,^F��\G�ͲcL�!���%�W׽Gg����ΥGg�w>�ְp1�x<:+���=��w?0����
<���ch?hh�[_��
������uXT  ��OH�����c��Јz�]���k��|��O��7ʈ��8Ѕ��i4��I_���"�)�e��+�u�����:��)XL>��{Ɋc�����!U�|2��4撚���z���l��1�;�O���f^�`g|�o�zf��M���`p��ԭie8p��מ�ץjfN�|�����f[��_��Yq��3��D�,�C�q�y���h%�i�d���PܷRn�1�G�&H�1f˶bT��j��1c�Ƨ�%�謭�_�K�--��]��sv�p�lN �.]���e,[���3;��i��.bc��hʜ���Mk��l���ǛI���j�'�}��$�Bf�Y����AE�ÑE`\�t�\�L���Ƣ��l�����oZ?5f�z��0��)��B�(��P}����s��z�y>��_9�oe����@���mT<g�n��}�-W�~��I��"!�}���T^����%�C�s���|]��e��c�W�L��o�E?�i���24!E��躊]�6���j�#�z��N���3y��?N��9!��uQm���=��?9Α�D�6��\���L*vu�
��}"�p�W��4 6��&a���A�+M�����p��϶��WRg�u�u���s��:��F#��ʆ��"6�hVWkZ�����������ﺰ9�rf&i|�%���>|��;r��b�0zb6-=HH��,�)�|���i��F�W��Y��K��������֓���G�P\&p�.�_�4��i ���IJ�yR��Q�C�S4���I�G��E�zu��y�/�52{��!C�:�R��\��{.`N��P[i)�}��j++�tC6�/V�Q9��z�	-� y��LHK�C��K]C�^���n�54!q,&�$���.2�s}�����&�CE���mY[EZ߿t����O}�*�2,!1������X�6�j��4x��юBßWǉD�CY�T�w���7�T��O��6�%T"�%�_0d`Y�0
Q"���4��-7Ku�9W�XN�7�Ǆ�a1��4���u��ᣃu��z� �_7�1xC=NusC��B�K�V�'A;�"�ݬ������N�	��;d�+g"o:�E����c�W��k�j�l:�WU�	�f�c�p���>E������.��'�u���@�����+���N�'��g��[>C:]e��A��Nk�������ݼ[��j�쥑H�HT>���#�4FG6���(�9<´d�Ƶnƫ<g��L^����IuQ �q��?� �'�3��bd9u"��	ܶi�a sr{�>m�Y�� T_�v[!lW�H���
ڗ�wBZ({�}��M�.&8,m^?IꀩUPj!88���%(J_��KW�`��$⻑R�y:S��Ox�,#�`�+���	�a�\1v��1����<<&��k) &��ln������W8�s��F>a�4�Z>s�����{�;���q�����
e"���6���P��%Q`9S���E��b�d���K)�st5�l��ZZ	����}u�P3@�tAQ��ƽ��/ys��Y�Ј��[&h���:�<��2�h*qq������E~,kDs��F�{8�U
���+ꆟ0��
JfU��oF���N����W�Y	JSú������ڀ��k���k���{ͧ�35C�C[�7��;���|%�Z1�u���}��Z�S�q�A��$o~���[����wsl��e�����p�[ם=�,���ī%[�d7��������	��oIc��U�+Q}Z⊜xZ)�6�ݴ}���sk���_Ύ4�m��ˊ��'���ʮ��'�eEz���!��M_k���@�RԻ�I�s����Y6yCJ4��vAπ6%�Y_��0���Ɍ����[�6���I���H���q�/�ӛS�#���9]�S���ݷ7�����e��͕n�_|=}���9����4�s;+|��+�?v�N�t<9�����=	{%#s<
�Kz�H���7���x�w9J���Ρ�7N�)�
��z/^z���N������P�v>_N��!�TqLj. 3�����T���<�Skl��.5�J�?�&��N��o�y�x�Ni5���}95P.��7���E����s/]{K��`���h�s�������W��<��Q�d��:�^x�Jq�ؗA���{p�?<u���܃�$ޭb��>a�37e�x�^��;��?�s^�c!���g�C�wH������ꨬwR�%����¯&`<{����b@�BDNb/���:�p�Y��B'D�)3m^S,g�ӗ��0��O8��6`b޿�`_�Fc�
s���+Ċ��4hY�Wvj�%Ӽ�aZW��A(06u���(k`,;�q}@��2NJ ����$h��<S�|R��By�|l�(X����(�M�Ҷkp��b�D��t��[�+6L��BL.S' 3�����c?�.� �ɞ!WS�4�IK�w7�����P:�ͣ`	�I��u����a���!��m>_����?١�0�.�+
E��ɹ���_�(c�0xP6�����ٜ�c?'�ã-P��⾯b3~��[��;t�o���	_�4	�j5M�|����^��	�~�79m�6/Z�S�K����-X���u��~�z�ꥋ�蹕��}�֕!�+��{����D����E͙l�{Sx����-��I��� ��<��e��_=M���ާ�^�5znY��k)B3�(����H���2\"_�֍�q�A�q���S"�I�����ԉ&�!'�:��zǼ�+����ȁ7I�_~��,;�n-6l���m�*��0����l �)H�:��c�~�>�R�Z07
v?�o��K���� �|mS?���>;�؛���������D��.�e[LW���C_��-�&/p����б/lҴn���l��v�����m���;`��Ò&j�+����B���9Čd��i�*��$BX��#,XR�%���~�����C�g�78y��g!�j��a��8v�4<f94t���m)�e̟�.���b>x텛�z����n)�t0�<7��!����CD0tqܔeVDu��Xo}����zT�U��3��=�6f�\h&lo�c&�rh�̷=�(�Sٟ���Qӟ�lΝ���u(^�\��l�za��#���������AFO'L*2S7`��U�2��8�H-4��N\VNpf�\���Gq�����VU�5(t���2���S㪠7�S<����'�^�v#��<Q����=0���w�x�v5����:�Af�����T����OFԴ�2��9���cK��U�5J�M�, Uv:��Hfz��у'STU��3��6.Rl�w��P�\3p��e?����7���>�C����a��[�[��_f�����\^����\��d�<,}<���\�,&%ǳq7*f�!�~�W�p�nz2��	�&7�)UM!�ϐ��O�g��U"|կŏؙ*i`�g\PB��e����:C}ʸ[��q	@�($��m)2c�VE��ƕ�s��EWPY��t�]��
�ɭ,��>�Fb�w������E���],N�ȃ���K��sl(��(�^7��j�GZe�s���ǖ�p3�E6��r:�r���V��K�IXu&����AM�N�;����0�2�.�5��~��ΨD޳)��j��;}_3�^n�m/�h±���gxzW���/����X�
��c�{��0��#KכG�3/q�l0I�i�(Jg��h���oLH���+:(|�Hl��csz��Uv�M]�7���)ѷ�r���J��He2�b���~�<�j!��U1MR|]�(y(��e���C��_
J�k� ��=�J�ׅ�5��<ho����v�R�D��S_�Z�3n1�|F��)���Xv���c��h��+��D�/!т�pv��Tl-�,�0��5�$tJUz��R$�$�[t�x����nV%��gp�ӄ�[a}a���)iD�ix�[��O,�C'=[|�*��7Qg�?�[PHT���FЦ��ӯU�B�\���"W�D��A�˟�4��*N�H������O�5��ԯ�/(����;ȃ�c^45�uU����i
�G̣��|�62�')����rɁ�R�U�D��f+�S��'�iN���S���9�6�
�U����Ü:{���梊^���\�N����c��+�{ڄ�39[���a�w��p&�ƛ�W��T�)�\�6�:��H0\!�|�)�ߚ��^!�>�'!����P,G	5
�3��j.���M6�}%u&�?'1�����ց��wf��h"�p�	���)x#���b�ۑ�é���5W��Z��U=R�:(���d`
Z؋H�+��2����@��U�dI��dBЌ�i��(�6����U�XW��J٣o����V�z�<d���LQ�wsTY��6�`7P�'m�m���^�M8!�9ܠ'.��:��b����;����\�p�zyj��d��dj;,Ƴ�M�!i�(b0��z �;W��d���f`�M�]e����@�E+�7��5K��������'/�#�����%�3�U�=�=�<�R�}���z�;�;���\�Ŧ�"���ۉ���Jh:�q���P
v��k�k# ��B���=�b��_m�(}����וG'���:p�p�Ǝ'?�z�,N��!��Ґ�xYq�ZC�}o�ڷ�h�K��Q�s��&�ƈp�B�{���eR���\��1S��l�xu�����+~���n$ns�����G�fbUp�?;.�Nz�(:9�?4��_�����	��4~�Yt/���s���E����3��x�[�ܔ_s'|�)��ʒ|Qd��+�>�U�99��mJ{���4��d>�A�Ţ܄�1B��p��(�*�Ke�N�4�m\
ܧ���D�i׷h��)w�M��'��{!(6\���j4V�M�`�+��j,�0��>�ەPm� ��E� ��B�g'ś�ޥ�Zv��:]�������K2�x9	�I��hC���(����m�u�a<3L`���xu�t����/0L�x��Ϣ�=�H��n�Kp?mIxV�u3T�6[,	�]C�j�g�ڴ=>A��'��>73�m��r� �������ns2������>ǌ��sM�|~}�W�w��j
�2#.�>Ձ�����2��ߢy��v�.��Ć�B_lu�.(DP ���\�vF41���u�?n�3�<^E�.^��W�9�a_fu�}p�c�o�O��z2E#�3q�rq$G���m�Km��4�+��o'�2���������<�:]�q玼�\�3ݛ���6���dU礆IBf�Rg,�j�+����@�.2� z1 ͚��7�ҩ���24�\	�6e*J䧦��rK-�/C8\ʢ?>d֧������S�p�ὤD)Ҡ��� �;�tiS����8r��l����]4NmU�9Kh��A]e�rE�U�lT(���L�<Ҳ��������I�8 �0�XW,����}�B F�p^�� ��9�Jfv�{�O��{�=J�7�r"���^}L�A�`AA1x(p�p!�u��/�����!å@��yS�Q�'�k��MB�M���R���|�>t�Y�ӬQ9��0VR�h����te$�s"�wQ����T�9���ʽ���օ
�9�a����F�$fB��@��O��r&'GZ�,���:##��p�������b	�Au��+���K*q~5�'7Ilq\�nPd�Ԉ����,��y�C�.2��נѬ��!L��u£�v��Ȳ�M����}<Yy-i��I�+��lJ�׬O}w%�e'��������I��ӕ�ii�>�.�+��ʀ��R���zE���RgJ�2�
T/7A�z�:���i��\NY�7�0�
P_W��D5ˬ�^��V����R����%�
��b��Bnq��y�����6G�|(I|���`f���G�,E��u��n�ǚ[����� ��$V����U��8��v����i��Ċʟ�j��re��}Y��t�O~O��Jn�2[�Ӊ�򊻖K��$j;��=��[��{Ԛɰ�:�I-6�qЅ:���P#�,ƃ͂��3����t=2��	n�DA�!c�{Lvy.�?����C��&��$C& �|�)n�c�u�џ��b�ՕlM�|aMz�M�+D%���n��6�N�9���3:��>O*�j6_~<UBi��*�w�X̟7�wL�Mji�6��{^��7&�v���M&�n�\ G�\�ˇRYm%�P�PP
ۻ�UCa�4�9�:e�iW�4	qX����ㇼ��:�E����:>��~�ڵr���ʳ�A�)*���\�/,��'��&:���Ý�4�ӌg��@F����e=���D�./���t:.�:q�*?	m��;O��ҥ7��q|�a����"��ҡ������:CÅz)���V��%1l���-|��D;;d
}��H�.�u���!��[WN�ӌ��3��Sl��=L ⫤ f�H��,�cn� AA�k���m2i�˞��_��8�9�h���Iڊ/���Tl�x8� �ߑ6�]�W)��h��+�e��7W��!�8a�VΚcN��h�[�w��AJP�,IzhV9�gt&�6ix��M}a�*P�φ���^�����Ь�@��7�R�uӴҫ%+�_����G��(��]�6Wg���}�LRx67#�M��%���TE���� Y�ݳ�_g+�.��u`N���W�oq�ş�L���U[���䋶���xGx�#�s�l����$s����5K�.Y�K�l�]=�I%&5kC#F�C(4�_9��f�q�@Ȫ'��E:���D&����O���_�R�����7��j��8."��?r�8bv¦�n�%�*K�b�3O�qE�ި�:��*Wz^����ox�������}�QN�@y�!�2���	J
�ߔ:��'쌃W^�~��!��,���ә3;w�2fW�~"�7m^m����r�A���Ksы:���g��'=u���>x��걖xe#f�����X���' q�����.�΋��T�M�U�ﵝ�
��Aa] ���R&� J��"�,y�_:�uJi^�p=���;��2uP�%P�O�ٰ�8�4ֽ�􊙬�@=�4Iv-������_�6iA�͝�+⃺�MR4T
�t�,!7^M��r��y�\wǭ���%xY���jLR��J[M�����(�?zP��*�2x��>zr�fD.�3��ZxF�?6�OQ�m�j�L� ��(Է���.���}�0��B���6.��t
�B=�,l�W���>� e��E�u�e���-n$��%�U���o�����l�֣�����c���H)ϷA���w��2;�Z�[���K�T9s����ҿPR�H�
Xx�3gq�E�'VW��n�D���4�t�{[c���wW�0����s����>�$�4��0sq�"�QHf��/����^c}�4���Z�=���d��v��z�tk�W��5V��~<-�V76>�x�����9J���~�z{�$�5�����g�'c
���OmS�E��u����Pû|�!pp�<T�BH[� ��'ܸ���a��L�#(����oe����-t��s�u
� Ri��������%���C������SJ۪^��� uN�ou��C[�D��뿻���i��M�X��4��+��]90��H�Cl�N
�M�:�]�#�ߴ+q���$��7k�Ft*����D�SԄ�}���y^��,"��JZ����ُ�A).�2C�{�Μ��5��K��J���,'8��v���uj}�'Zq�HZ��\e�	�=WH�@O�,mop+W�$�q����}�������Q�w3Z-�5O�'�.֤g*ӋΖ�sx��q
�n��1	�[:SW�y�yE5�Ԉ���ǣ��'y2������î'�cV��Ԉ_ڻ,[�q2���+�7��g�$��++Y����|��3��*9�TʕFS`��/�EwWT�̌f�:E�}�������㽮Y*yf�v��CW�@}��\�@���& o�Ĥ ��%YrR���ѱ����xM�	��"�$�������f���s(��t�� �+t'rí����=����Wv��I`��Y�x������yxqG�p��Y�6�u˾F�{��<�˫8E�]ǭ�5����4�A�F��W5ţ��������r1�wk��SG��ԁ^���q'O�BM��gNOHvm�A��SJ�(~��|�_�A�G�Nþ��N��Y螌zG�q<���s>0����;�s��N��\�w_�W;�(+�K����z��Vd�?Ӣ4�§di�߮�,�ܕ��&��v�3:�͠�%�X�d���C�39A'Y�CcK`.C��y��#l���w��`.�~<�Cu�*�-8��Q[2݃���
��GD��>tr��~Җ��5���o�T>��`�O�k6-��zbSZ�4�ӏ�-�i��K��X[&i�T�e���kЛ�3F���'o^��*O^Ɔ�8���o�w����|�Y;�J)*vp�ZH���s;N��?̧X��W�=�E*:��7;?F��M�ɋ'���穅���un3�$aK����CDCjP��3�L �����/D@��ˈ��_��se26�jhZ-k�R���Բ-&�����o��\ ���t����H��4B���5��z�W�r� [H),��IQ/�c${��D�/`�F�jԢ�Ey��)kR;�<'��9_:9m9�+��|��,�)y��װ�� j���X_��o=���r�o��9ϰf�Z�Rԁ�� �0~Z��>dFX�;�BH���
����gְ'qY�C��p���+0I�m"!ů�<�<W�N|`IO�#9�R7;l�Q��<dx.����+��.B�tX��)�^�Q(�-�Ϩ�<�$� �3�����x���,�jZN~WͲ˻X��;�����c�<���j [!coSN�Kk�c�_��KX�]�ZJ̯�G��S��ڽo�8y��+ek#�8`���p�q����-%R��tI��m~�$�rq!NMYa��(���I�b%%��H����ܾ�����<����@x8Y?�O[�p�Jr�
�bܖW<%�|뛓��"�y`4/2��9[�lITo��Q���w3�k��l(v״t��:J7B�x�5������8�= �d�umn@l�������h�Pԥ����� ��J��p26���u�]J�	75�O\|������y�\=zY�4l7l<�|��~�&�n�&B���0G	+���Twǐ}^-�f�`�sT~��Co�/0�_�\26��ܝC��⢑lB��X⼩�=�;�ψ�S�;��b�y�C/.%j�u��h�][�w~T��`o,]��\ 3��F,��������%Թ��%�m�>�,.�&*ԧ��%���=I���I�ۉ�f�7��L��s1���lJt�&�/���R��+X�G!i�]G�	g�F��2���ANvv�^����9/�,'�l��Ff�4�<-r�k8R�8|����D�2��R���P�Y/��]{uu6���6��hx��n6SU]ڮ�~Ï���> ���^���r��,��%x�E�Lm.��m5[reO�rd�Y>���y���A^\KC���a`Y>�n��b�|�_��^�^��nЕsA��b�i�]%�)R���
-	RX	���p�.LǘDS5����;D1՟6�� �c�=F�Gò����죴x�xѣu�MGOə� u�pT���̝�i���U�n6��c��$�_kȋ�ׅ�\�W�su5��d	���qrԘ�l���yUsG�*���!��D{{T8 b͌!Q=(n1Z n����_�����:�Y��W[��'����(O����5����)������!�6��>�w/֎���Ȩ�;V��~-R\��}���\��M�J2ɳ�a�j��M�y���c�9���j]���+�-��";�q��a�l�{SX�7�6��4���:F�3aj)?)�R~s������_�&4���~�^f�"�Q	�..����u���'m�Р����¨e�
���3֪��9�6G*�j�U�<�?����%�ja�h4��O�2|o �;�E��9����8,�`��D�wIP�=,�+�I�w�����+|���8p�i�J�o-ԓ�e+��rde��I!1��hw�.��A������{z�PrYjR$��͸� f�I����`w�ȐK| ����EGs1����!�)8�BU5�4�&�gc�0+ �?����X�ߒ{I��F�ƴ���l��ZoZR���ޅ-���>��!���׭��g��3Ύ����"R>�� O��h9�I>Wa�Dv Fi"�<�p��AsW;����R�k���gh�R�N��~0I:W��DL��0.L��%��g\T3�b��C������U���A0�����Ckw�|4���oӿ�.jۍ�t�%�X0:߷���zm5�&S�} 	�����V�&a�����Yh\۰�k`�2����f"W�^nY#��|���8�KI]r׬���7���y<��#cW9�TY�tH������&z�?M˝����������9��NO��/V��N�J�w6'2���~�"�\� ���X��:�#J��'
W-�*�/�O/K���|�#ؔ�
TlR�fT���p����3eP#c�~G�N��W�E���f��$���NO*�52�,�O����am�CW%Fj-p�(�3}�������HI���  ����co{�Q�U�?Q�^"Â�zL�����T�^-t�)%�3��D��uE�ѩ.l����2t
�<�c���:\�!R R6(�����-���$�&RW|T�Ǫ�A^���7�bbxM ��������l��m�n3_�|�;ګ�y>H;�aF��>T�ER
��՛���g�b �[��:�GAZ�Eq��v?}U쨚�P>����ok̟��j�m��N.y��@��f���ÿ\��*���!|�7~ԥ̘���X1�4�"�������覗�EM0L��B�mg�	W}Hf�O�yl���e[�����4wYl�_�^��MN<�WŅdj]t�u�e�C��׀e��EYT����I��d�sd��ɽ��8�z�c��SF*�DM]��H�F\y3�(K+(� %�_A�@����LJ����
��`��o^m����d�^%�¼h��22��LW2�|ɴWbI�rZ$�����qGG�d^���h���"hjdy*�5�w�O�u�G�u�b��T}T�*YJ�e
l^�ޥ�Ȋ
���'#�^�3j�hF��<b���p_OA��.��?�Rϫ��s�)�B�Jz�R F�-9*�(Zt@~���yb{���0���4tp=6}-6�h|2Fp ��=)Nz�Vi�m;<?�8 �L�b�p�rP�C�A��f�LPs:�v�G�y�GS�%U���j������9'�ANi9 �4q�����q�a(�3�����"<h���g�����I���]����K������a����n��}Te��z��͍���C§�?V��F'K8K��Z�G�?hfҲv�jd�,��v��P7A�`�f!�V]&��Bz�H<S?��\ꥸ�����,"���MW6_@Wv�������/���F��
�3&O�(����,t>M�3wV�{�2d�oŧF.�&������"�,�+�m^�*K�},��w�Dl���[���v�}�nU�(F�Cz4������3����9����Ξ0.݇&����}�$��?�+�acN~���I-Z���4��mD���L�=n2�X�w�q��-�Q]HU�f��\��-��ҽ�g,�XBM���^0�9��f;|¬0�8/��߉���oïr|O�
����������~/,H��Iy��n���(���5�
�b4����È���Fp�H�E��b9�`��a��%��R�����.2~'���mj΍���c���y)}`��./
�0j���e?1�3����5��#�Eư4>84������7C?���p% 羑��*�v_���0�J���ԁ�+ú��T�$�a�d��4x�B�Mv��Mu�.��I�R�.���#D��/�̕����x16BX����C�8�s�Ŕ[�B�.;�^�BF�oEL�A��
�7>"Xynˋ	��x��m�z���P�5��� �P]8gP��;�ٯ�F�I7
9�����i��(�^�
3�#q�b%�ce=�ʦ��e���p���Yȥ��+3~3w��� �Ek��e���r1"C�"�A,���P}}�3�Ƴ���?ȇ����uuHh�Mjs��K1��:�:�6Q��-��D��bx��h(J_}��U��>�y��Fp�����f��S�*��e�9�DJ���9=�lj�X!q��P_�\���QYSŞ�)�V\�����-G�ݝZv|%���P A D�-���� c��H�I#���� �|g؞��T��r�.���d�z/#�3�ʂ�K������ķ�"�'΂dn"�X���P{�`�ы�7v�Jn�(���2Ԟ0=.~s��D�}v��E�=�r���X?�}�3{G��o-;�
s�-���]r���$N7J|%�8���⮲�sok]�&j�J��Qp�s�Л�
�L���*\"��f]@���ME_+�;�6���^(��I�/�p$�[���/�%OҔGG�����D�����ڢ��{�?�*$�{���ޯ���',���F	M|���!eh�v��������X�(ȝ�O���M~!SeC)���޴���u�m���_��5��?S/$+d�ľQ�Υ`�+
0U��� JC�0�W��l��~�(dy�}9�B,0�8[�쥖��0��B�?�������"d�`��~F�����i�M\����?g�8��aa���i�*.J]���2x&�����ᥭ5�y�NzE��
@��v�,(C��?zn��9��K/�����}9A�S`:�9�܄���V�*D�I����xQ�-i���fP�	W� �+��)�|��V%������_�6� �9�>���=�=�II^���'?쬐��2(�Z�{�-�����˰1W^�)b)>����z�����˶e�W�D!��f��+�,�]�ǅ��>�|�iIS���2�������JN�<�����3&sU�g��Kb�{��W�
k����6�xH	
��͝��
+�t06"�,bBsݖ����Z�ֆg����M��?�"�(,j��L�O@ÕGI��QXPN
~r5&�l]h���-[-������;���Z@��Gh�/
���b�f�`bg�2�'�@���M���_����ZI# Qt��<�Mk))�a172)��h��������D\��b?���n�V[��3_q_��ql��=jЌ��y<˖��B���0j$-���bF��=iȺP�jkX�LAȒBB._�%����#/���o�>6��+��bu�ƞ��	RI�}IDO��h�Tb��%p5�y��^ ���s�e�yu��_x�<�+��$%��Խ�wbq2��H������G�bcu2�R���9OP8Y�������Cܡ����*�/Ws�W��XZ�Њ�yX���rW�0�&�t7[�WJM��<��!Ï.��W�~�Wz#�%%td�[ۆ��\�\/V��F/���Z�WyK�Nǋ�wY
�=w�>�X#��m���<:���C�F��W'B��`蒍�k�Ms�Z���<J�+�s��]�
�p�I�`.`�# I�y�֔^��%�>i>�m?��M��7��z��eђ�5�@��A����c��@�+kfF���P蕖_x���m�֢�q��/�4cN�ax����!~W��F��D�q-�o@���� �$Jy�r!;	�97�;1w�u-�R\M�A���PQ����qQ��3H�D��[CQRvUh�.p�,�}S��5��'��u�PiY[���'�= �УdН��p*R�����=�5f�aɆ�CGG�Մ,�C����c!���t)�������H���>�<��ħ��C���U\� N�T\�%�HiLB�E����� ��~�����c�<��Jda~�`0j,�B����~#4�q�4�M�������.!�=��k� V0C��JB�������+@���@u^i
�,�RɄ�p�*�f���sC�t�Б�JW��	$E/k��!- r\X^^~�q
#5u�f�˨1��ʧ%�p��̣6*���YZ��E�G�$O��ēs_N/V�����Bg)tޅn�$�o�^������fb�Q[p�&�pg�E@i_��X.�	�`u+����5��C0�O��dDS�T@�f��Z�R�>5��V��T�>��`�i��ۆ�NB��Ǖ����Ч-�3S��e�f0s����\ﳉ�/�<�JҼg��ij|�m�[�q�=�S;�jI!~�9�X�L!bv𬶚�5Qu@s�|��0��\�Ҿ��b�s�͈�ς�lw&��)� X�iG?�T\`\gÉ_��������}Á߫�!��b[*@��9�`�g���_������nG���*uR�g_}�_�l��|���|�.�^+��&S�a���f	�!1o�#�܉�:XcY:����_����t�_�R8rqF��O��$5�+L�<�����P�{q����/f�ʨJ�h��J�I����H�(�Q&FVq����#���ò(��g��~u��I�@��8�v~�2fG�hc+=�����v!���4�`�͊YB͊�]`�&ƾ���c�u<��-	�Z/;�-#�A���COb��-���	���Y�<J|ůq&-8SM���ɻ�Op�M�PQ�=��Iܕ� ���ϕ��+�Dyp"a�ƨ-9-��4�n������� �Ӥ���wF��y���QR,޼o4ͣ��i�xs���Y��Vt�/��/���>�2��E��
��?p���^>���m�ן�����̾��\d\YEwbҌ3x��Aj��f���OĐ��_&�6�f�J?BX9.�j�Y0o�)=�1Lbh���t��\;
��|�'�DvIF1g�xQ��tꪞ��H�`@�)��w�����Qm��H����M��옮YDi\������/D	h9��^��lG��Iw��\��B���I����r�)�6r�{��O"�i�_�ț�d�ZF�я�^	�����]Th���4���t6�!8�<�ý�1��_`��&�Ӌ�r��yK�~K���,s����0�� �Zo�|����F���ۺh�ݜ�ik�ä�7)����ɘq�&n���Uۘ�ոg!,h?��{e-�͓d���i.aC5XF��N�)�[.��?���p���7�GCN�����LO���kK~:�/,��/�H�ѣ�4Y�jG��0Mޠ�F�K�7�KqA���%�D�0sH��h!��X��%�,o����d��o��8����-!�e�8'��F&[�^!Ό�ʘ H�o��b��U��X0�cIȐ��J
���R���������1�!��J�,D��S���_G	/���E-f �'j�ڙ��+����i�j]Ɨ�eG���W`��-�&�X�r�������V�-re����T ��x�W|�+}p���d$-!�-V��#<�g��b�x��	B=.��}�n�����?�-Q�2�I<����%49(�m.���P�b=�x�@����n�W5��|��|��4�"i�y
�.Y�v!bX0�M�|��F4]�����ܛ�ZI>�����Ӱ<-�{��#�C_�q���>ѯ�����bb����e�U�$��P��-�����ܜ�#���`_�&�e=g�QQ�E�ץ =�u<i�mK&[���4x��9-��xv��j���B/�rYS�\��rsw�� .k9����.�m�M�ɑ"�D#'��C���yY]�\b�����,$_�8}���$�\�������\eS�EB@@�P��$��Z	i�f鎥Y��nX�Eji$�X:�i%����ޯx���tf�ܙ{Μ���qI��f�u�|LO�Lb��`*oG ��@$���w2��
v����|U�N*��;��u6�w��U��Y&��[_�#R����I�SN��sq��٨f��˕M����`v����Xa#O�w�F���# q/;��2�_����A����&��Z&/?�K��`Η�)��u�f���'��n���Ӭ�����7����0n^F�L���vߵ������q�]-�V_43��i�^����cxŕtR�NK"�r�}En1x�+�'v���.�ձ�WW��߸l�W|^y�J�>[I�!�Z�0�[tf~IW,R��3���N��Z���:`��QB��}�0 '`S}<Ks|�5�dZ-�����*����b*�{���,4��p���~:���[P��bᴸ��i}��X¹qc�6�زw��.� �--ި��<,ۉ����ڜ3i�`��J�f�q�k�*��T5Ê�w\CaE�&�!�=�ا��Ob'�cv�87�$G0��4��/��N��ȂEq'������Y�?f<��'i�d˱��Vt�i�p(�|-y_T�u�vf���h������gZgn`��4��Ҳ���:Q��}C)����U#��uE\vdoWD[���j�}vE��C�R�)3� ��y<nx�:����#��Lt�֮+�X�l�f��QI�E�L��*}���-��Z��b@Xo�F���T���GjT��Lw��͇Ad�����Ƣ�a� Љ<I��k����[�q�va&���K����w�S��V�o	��{���|{�@��AZ�����M�W�M�:��y�I�@ff��h��B)t�W��t�CH�Y��1M5��X�,)�7�?��hCIi�C7�,�� ˩Ps <&/��%��)&�+0k¸���k<�[&{0��+�1ܕ�$~j^����E�U��c�"�d�Q��R��F6#�|�8��x,t6l��L	&�W�,=���d˨�"�J���%���vCCRu2I�|�s�ӽ�s�EB�e#�� �O!T��z��(ߏ�K��Y�!;ʟ=�B���R����6T�24#ݲ��2�Z�(/�Kķ�r:�6��Ĭ6}���"�,�ɴ��C��|)���w8O��6�r=�HM�cVvv�{	��̝��p��x&����Wۄ�8&U	���0�-v�K��W�aVde�q�V�ع�T�J�2����#�2sT8�� �R #��E{7M��G�ީ��4��;���}�HO	L�3���	tW�9�_��yR��њ+q��\6�Q��)7X�(�j��?}b&��{�������n�p�;�~*B�-��T�I,��x\R�!�w��WL�Ul��M �Pa�}�������h�91QӚ��SMP1My�\X�C,z>x�2�΀������ġo�g�F�T'�R����[�U�4q�,����W���n��d�릻�Ջ#?�S@�A�<܌��)/��ƿ	���|�q ��Ҷ�Ͻ�_���L�,ϴ�Qh�i��D��RQ������P�{B��W�K���b���8q�u�I~{{�z��J�ı����2�)&�!x��E�H�"rǗ�;�l�YhT6�E9��;�{S__e+cDM�Zk��i砙e?�JT��ʝms�Y;m����,�F�c�Ea1� ���]w�)�P�A����U�X
	�Q�$�鳌�e� �<�v�[	�������Y�_�㳺��i�5Ng���C���K ����ջo���K�[��X��"@�:��D+F]|
b�~��h�=t�Z�GPKɸ�PA�O�����ԓ�����N���#~�3�sFK�-��F���HP�v���tx���x!� ��j~����f��jԇ��YD+�+gZb&��|�yk�Cz�Þ�?���}�?��S�%�1��B�x�)���<�q��Hw}��K��[���j�e�J|Ә]¯���]�޲I&�N�z���m*̗#�%b
O~�\�X�ͨ :SE%zZK+��~��[]B��H?�q��?F���e_=���a{D��cF'���1��y}����[O�:�2O�?����5��p���ܽ��jw��"K�նĻ5����y�{��̉�@]�6���.�A_d�BYB��?u���%����'UO�,x�$�8֕bۮW�@n�)iׅF��q�����I�^m�����s�VTd�)'Ֆ�$f|����v@�|�J#��dŻ7� ��ɯa����Nw��u�0��u��|n��&u�q�7 �Qt�MY}s��6���]�`z2���d�	�s���9	��]?c�`�6�_���$P&��+�D܃a�T>mc���1I��ݚ/�׷ش)u��xO"�����O|����a{{��x����.r���J0����*ň{�S���h�����귻�p�Ad�ҜT���[ U�<?p�� �Lf4س%~
;��yw��b�őy	�C"��;��P��\�v�e�C�[w{�<p��u0n�j':�t�ً��e�/�T�)���|�#w;m0wyF�j` �6��@=�,#�|XꁾViq��n�"�Z^��C/���O���YjT�;�z��W��0�q]��lUj��8��%��3�]\�ݙ_�^+tϔ#�f���.�;��=����`U&�d���b���`bٰ�9�}>ۓ��-��.�h�O����"Xy��d*P��3�2.?�����������7`�?���ro���nQ��QS��fX	[�X#.:
qTU�!���<�e/O�e����LQ,\.���T�Mij�݅ѿ�X�׶u\6���q*zTZ,�0��ql/�یߩI�+��#ޏ�}�
�
�ޏ���h����������E류�H��~j�.W�y7�����g[O��35�a�=��-%���cK���p^�j�����wVG||ў��6z$czL��p�N�*E��d���8B����2��[��*���8��NO�o�6���~��%m�;4��^#m΄��Ph�0~���mIO?��m2�:h9L
�d��V�F+z*{a~�<�`%�	L&�:�r 
�gO�4ex˶NHP�_���~��9����ۇ[q�����&Z���(�%�?^��	�z�O��(Ґ_8H����w]^=$��Z��F�?�[zl�?�p\��}'h�T�c�+"�r�H����>���S��D�NZ���W>v�$hς_�� ��⣙T�̓ͱ*b".�@�����Y�a�I�Y�CQ�[�]�~����3�7�g����'8Q/�,C�=�$[��+�b-N�%ٷ�p�pi@\���5+dD3\��7R�3X��BQ��rRd���X0��z?7%ph?�*E��L�5�i�x�ڎ�	Y?e`�x��]��42����i�Fsk���{���탞�9��T@跦��޼4��������������zm��=��d��6��ݬ�P
A=Q�GL J!�7�����Q���j��� ��vf�*���퐅qi@���/��FD'����ݙbOc���p�����y�ک�J�h*s-��9����V�zu	�T ��hL�Il�0X!�ME���s��%wm��f�n;OJ��,J��9d!�8!�O�4�F�N��ׁ�1�s���&�@L��ہboL\��d����a����������&�u#I����Q�Q8��l{�r��jC�P��3���X�z���B��*�����H���:�F�M�A���MA��{@E����ܘ�Y�-�C.�2`��5�/��~!�g����0n$�o�?p'0�fo4<���!�H�/o�pći՛ϔ�0V0	���jU��(U���-lS0�c���%gt����8W��8Z�����aM8,}>�hX����Ӓ���է�/���?�E�1nL��=Wң�,�.W%c�PK   g�~S��RC�c  q  /   images/e1605cfb-dd4b-4fdf-9f1a-7191204fc245.pngd|uX�A߮�")(%K#��� ,�%!H�(! �,���Һ������ݝ������s��u���/�P�>έ[���_ʨݺ��u�v&�V~�N��.jrR����Voݢ�%/�\��hc���I�Y!><�07ջ����墳N{wD�n׍T�77�����n�=�FL�-�lB�i��}Jا0�����E.�h��V��kq���í�t�nc=����h��O\�N�>N�<��/�-�w����B2��c`�os����'��d�p�Ф�WXzfdfF4��
BJ��<�Dݷ�p�8C�ߍ�����Χv�B=�,��<7���Q� �����VmG������>���y𜧑�P�����X�4�R�t������hOz����4~��m���.ɉ�2̇�f�07�ܣ�?����Xnm�����p䫓��]�3 |iD��ҙ�*^�R�^�wyFSb�X>\s���Ͳ���d=Qi���ׇl���L�+��(湷⹿��c���J,Pg
첧�������b�οOz�l+�\�{�քzf����rBB����~�'LLL��)q���?�.˛��b>4�e�v
��=�\���f���'i��Z3���cw.���x��U�W�Q�:.��>�!V��D�6����W>�S��p����$�u����m%�o5�"1����~�?V2����+l���8WUg*���ɾʄ>���7����}��{����Z�}�U�"�:�ܺ�d�����bdd$B������Z�"/#s7($d���x�/Etw{�Q�Lp}hZ6�b�`oϹC��:)�Ə bbbKF��>
�z.++�Qe�i����XV���n9--�����d!��߽�6�+B��X4��"�=��i,��)4z�$	��t�N��H���{6Ym?���	�Tm,G|{4=�ms�<�Jx�%�'��_=��TmA��!���|��8>%$'�қ/��"����jx�B��,��n\��|�:PANQQ����<��Bݼ�����pI���o\��L|wb�4��tk S.����ߺ>]N��$�u)j	AW!�]5�A�O��|{DT��CA/P5X-��R�ņ�lz�ߞf�5R ��}?R�/ǮU���g�31~�*�a���D�'�%��(��J�!+ ��c�oWi.���+�[��m��9��\��J��,h�2U���X��w����H!�bo�q�T�(=}��TS`0�+�$1�C2|ӯq0��O����U:��r��)o[{;���`ɛ㭩b�Z�m�ct)��.ނ��߼�2�������x�������su���c||h�H��ozzQn7�[�Ϟ��t�݁�C	ѫ����-��6�XS�ɕ��:���&���~�?�3��ꈢ���srr�5���Z�bٵ�ޘ<��#�����ͪ]l��x�wJȭ�Ǐgkce�*�UJ	OMzbX�-,f���4���X�v�H����,�@\ L�wus�|�e�^'�󾛨T'�u`U.g.-��Yt�Բ)Y�*Pa�k���{~,��\g��+ �Ƹ$�F�M��=�C�D�(1*���5y�����>˾1V�M��g��J��H#[{{7%Xm7N�;>~����y�JNVv0���js����r��}�/�r��f�J������D�_�<��|Ϗ��������mT`菄^��O��z�Vs�v��%56T��{�=V$���G��l=��=�R���o��QЯXv�����X�9����	����  _��&�'"���^Eш�X~�̔F#1�oQ�����������i�oGO�'�}PI�^{KvE������w�G�����jU��8��]�6nz��WY|�o��!!!��%z����Ĥ*c�"�H~�����t/Pؽ8�,;�c�^����9����s����_��{h׽��(3��fē�t��@������%�i�G ���Oq�A��w��l����-((��_���?z���j.$�c����x����'/��C�ۍ|<�6��3)�x��G)@x�?� F�\^^��U<$~�N��QJ>�˄Z�:3�?~�nn~�y�/����w�L����Хb���\����&_���t����.�4��ڟ���6�L�����0��d���>��� _}�'��`e��,로I��ׯtN���7�;����mM�k{4�k��989ͦ�|m۝��BL7D�!�ҹ9Y�O®�(�wھ_�����*���L76z�7V�¯/����_�v�?2D��(��l=�t)	���E���Fq kQl�9���!���=i��:����`5��:���Џ.Rްg��D.S�F�s�+���$�p1qq>�k�l��b�L �j::cB�f$1r�E�q�������ˀn�̓�_���且��۷�--A���es����QQe
]���΋\�uo��z#�d��&C���p]��'?�����89��wD�*���u-��IΓ��?��uʴ���7�E�P��*V���I�)�%#3>�� Ać�t�-P��c�:�=�]�k-����@{� y���a��V2��/��??�u���1#5�*D�g��P)�!�mv\m�_�_\^��a��K?--�\�O4� !���B�P��˯�|B�\wШ��T��;<%e&��)��������5�3�u�v�G ��T����D�~��zB�˚��e�h�ɤ���)I%_xvp(c�I8v	�۹�Sҧt,�gá�f�^[[[R���7�\�뻍�J[XX�M�L]�>ٌ=��V����2�hsR�}b �
 Z� Xr�1�9��Fp��<�Wڍ;*f�i�Z��G��!;_"�!� ����(���N�s��b^��XDDD�q{1�@���� I�aG8!:[gƁD��ڎ@%[���ء����;��I�#��*6 �EC&.S3w��@$O1�	��}�v��t0�*��".k��Y���耟���f�^�M�����[�X>CЈ�5z-�D�#��W~�KkdȄj�M��*ఈ)��`(��G`��
C���"�ȝ�͕��'l��s1[ى�s�O*y�u�0Ƚ����K�Ԫ}5$�
�O�*�_� �� M�q���S�}`��*���5����W����?�|}*�R��11� �*��7�d��]4rn���Z��B��;�?E�=�g����5��ݎ6tG(ԋ�'*,	;a�͉.�<a��Yc�\m�δz%�ԗ-�~��l?�)�)ZW2���?rSl�}-d֎G!�V�\C�X������jydkk+����N���0�%�?GD(MTja�ۨY��^j��7���NK�����~�]����w�UN>�wV�N���Z:O�\.b��� )9���Ϩ����o�5���34t-��4���s�%ȩw�qӨ%q>C�,���������8]y=���Tȋ?��|��[��4\����ț�]x���5_����C�B��'��&J-�����Oչf~-��sB�&0��"R�$]c>��}�p�H���%�)'��nvܺ�5�.��p_������w�Q�׆�7�Y�5�x���e�՛��5�|�[�2dw[�\��]1�XPɎٛC.�V����/͔�U܇��i FM>����5@Y^���4�)�ƟB#�
] �P��%|N����5�ﲤ���3�����4TS�mh���� у~�A�Қ��ZVYxX��q�`X�C�UGxh藷v�}�Ľ�eT�8���a�����銱��.1�Lw6�I��7.�kQ�#�0y��+������������������� UU��W���]1>��/8�6q��G�����u�k(w�ᦙ�K�0H�8���_�1�%���M\�c�I���a�82�������W�e	��LZ��i����G�=��w��� ���#��͏/�Y̳v �#E�{@�� 74��⦼�e/���u��7ע�̴�N��肠 (���s��8�b�j���~��߿�5�}s���8��u�Rċ;hT����p$�&����D����TTT4�5�8u0�A�$��%��#�GO�s7�9Պ#q	��[�$�O���*
�m2�`��g��L���J�C���2~g?Qy�>RD�ֵY*�����S
&���G ���۠A>/Nj#��:��I���h'�X�W����B��%0�?efr�}�Ќ�GG��� <��m���Z�8����� ΃it�DS$M� <w��v�a�eh��Xl�r"~��� ��< �w�������XB
l;E)���VL@��P��Oi�����8��l�ff�t��EFrXr%�u8Xvׇj�J��\1���U6(V#�I$l��`]������^1�=ٖ�F������`��5�w3,ܘQ]��������5��W|�����De��O�����3=�q����jL�$� Ё}rr�ݲ�2����ac!�g�_7_㓬�{�@�S�;���ܑc�Hd�^���1>>�#����IO�ܣb�6$�-?�M���<��!�r�7$�D��(���C�a)�����5����ц.���n�a&�������1�2S}�,9Ի��L���/ ��3�)�����zd���E9QV^�⼹�V��S�["ʲ7ݤkk��:��BRD�N1ЗU�S��3�+������U��ܹs%��F�yD���2*�3�r�]�>��n�]_]�g��7�,j�FKf�#�DR�j�Y�&-g�xl��8���R����?���<01>�
�,��`�.����Z%"��d^��0b֌�*^E.�ݪp2�r���y���M���N_=�E�ޯ�gmM7&wtv�~Ѹ>;X���P����v�#Z��Xb�KK�H�ƺ��Տ����������Ņ�R�mw�R�l` ߙ��۬w��54���
����
#agѯ�C����K��z�U���N-e�i�1�N�|������o���̖�jb�"�̬�r��꺷�ۯ�h���6pݪ�C`�u���kk�c�>��%=�P�s�������:����A8��j�C����W�)"�V';H)a�-�
�	�9� y;�r`E�����Q�Y�B6�|V$Ӈܴ���h~��#�/P<R,EE�@��z�@\��F�c{��d3�I��j���f?߮/!�x������%�I��{�qpvh+ȣ�%����RЎNRR�~�����X ��@f�
�^�y�Jg��`��T�{��Ervy؊<�J�V�
�}2j��QD��t��6�{WC]�f�ߜ�TS����=;\_l+#���x�/æ4I_ $HV�z�#��A�������t�g>�R� 	Mś�AJuoη�ʤ�0,�������Ā��uw�3��r��бv��ь� �(���b�pp�)��Ƣ���'��f{� ��+�z�ﹶ� _��6c���GW��u~�nQWN� ���xX]ڥA!�ד*�������Tfq~��v/�_��g�/��.Cjۡ���e�I�Dm�_2dA�<e�*$4\���kR��[E�]�h�3�/�T~��_�^:��鏮���|�Ի�GZN���8Nv�gc�;;�|��!��R�1+� w)�y��������c�&�̩�
��
&i��sA��o}}�!p��$�8CK��A_[�~Ia$4�� .��r���yuf\���7��G� �c��U��I�	��  $�x*E�q���L���%j��3b�>��,� eix�$!G?��vWX�6!��'^C�K��BBBT\_��]��ZY}�	�\�$2���6�0�=��	�Z�?b�{�\�����A��3{���ZD�^�	�����|n�pv:h�����Fc�c���KߵHl���`�=tq��*/5+��g��k�R���x��������Dh��� ظƨ}Mr��W[��lA��f2N=�g6����Ϫ��t�z���l�����l�;��<���_,��#ب�JW3�R̸�A$T�h*'����ZJ��簋��~�"&f ~�{�#���b<&a7�2�)�v�?���]FFF�ή�T�q__�)�h�?�ƴH�鋤VP�=,	���i�0��������$,������Hq�n�樖Θ)���a��E/�N�R֔��DZ��n�����rİ�����L,P����60��l�n��v[� M�K_Jpp(&�o��IL*��F�	-
�>?D=\�]�0�K�����iVO���,c���&`���C䋨�o���
	����/��*���
�-�5��	/��+�w�L�4*�|���: ��g2�Gm7�l;J`�S�x������ż^�-�poU�%����xs�E��̱cX뜍:\������3�0��O�B�,���d��c��%g>\|-�S�/��Z�|�׆h�]׈��r	Ho�'�������y��OIg� SZi=�<�P�å]�}�x�|.�������M���|��DEۇ�#OI)�w�.c3�/�a���b�|P(8���t�z�iTnmn�?���˗/��]�x�� |)ߘ���d���%x)�������+��1"ob[�R��E|Q��^/y���570o�^�0wh����+|�?IU͸��^��������$���v8.)��1 &��O��gЊc��+���$��ť�P��@���:�K/�{���\W��ٹ����SS4o�ʊUc��͟o��t(9�_ʀipW�@�3(#�q�3�Rz�pv-�7w���l&*g�rL�hc�{cJ�N��WHZZzzfF2$3s�W��%zZ����v3M�Z A1c�?�e٠��Oj\�o�ŝ鸱�h���0l>r>��@��b��
-Z�zߕi�U�n��:���*f������r� g˃��*�1u�6���6�_����ͣ$�75]��,캦1 ��qDd�U�#�dD>j7��&�Q\�q�Ԅ����3J������S���oVc��^zu�������*icbo�D�d���:�c=[-QO��] ?K��99[=R d7�{�^�#��>	xg���`a��f2���/�����s�u��Fh��d4�&�z~��t�s�WX�6׬�D���9ˋg�PԖF�����u��D�yYE�g$Eakkku�:��wp�Y�ס��z�ůvD' Rbb��d׿�w��[ʿE�O?M��0ҏ���U��
H����^E��b��I��h�ۋ'�a�T0 v��.N3��O�Еć�6�������G��05��v�h|r�z�7�<���A@�6����)5�C��/�u��^����d�8�r�PEE1�0=�NOwOw3�
��=}���hx�	Ik�����]Q9��7<˻�lA��"ݎ4rp��ݱ�ǌ\\},L�ƞ�� [� �é_��J�E�$a���_;�vv�}ϏjQ�q�8?[���	0Z �n�2ϯ#����8�İ�n���bXտYTR^z B}������4���VX��'.KI��K20e��#W
�4��s���EUy�vJJ�u�'r)����F_��ȥ6�iu���y��?��/+Ȱ�B�x:�����^www?V���a]jv�4�P����] s�TӎaW:�K"��߃ e���Q�zivq�+yi>Ľ-A"~N��B4��NvL+�C1g�a�"f�h9V�s�?E�S��X��YF��"�t;^L�z����G����*��#�i�e�[��_&�]m��vke��!9�٬"=-'{����K񌌌o,
����jp�}y�z]#�$/ewQlX/����[S�r�����]�K&��G4����u?��/"|%���y�<'�28�z�u��9NV��Jۯ��oa�H^�Hs?}
��͵�i	!P���#�ȗɅ����4J_��} ���F�P����A=�P4x{��WVyr����!�][v���Bg���H��p�h�q�cn�\�<5~�-�|��	�f��UAEƼ�#�iF�2�����9:n�A n��L0!�шp/������S���pg :V�`U��~�
aM���AA�����Fbr�
q=��G�
���{�f��9�]y��2�4�%�����IJ�� E���t�����`�Y�i�,���p� �-N��D��'�˰�7�QY��TH����A��P���w%�YvE�#-��E����%*���o�L5�;�2Ls�[�7	�����uL���ʩW4�w�iW,;�C���z�K̉?ŠO��H��Ύ�5�wx���́�6��"2����L�8 / E��w�Q�-�B&��B0Xz�~��y� ��d��=Z>ol/z�VVNJ�'�ry?�O�_:����/������aQ��B?��r�R�v��/�	��;}H����%>Z����*�d�A�p��+�y� ݶ�e���,F�7�q�m�rn�ӗix~�_��[��XYz���*�B����?Q'U�K��n�<nM�.IO��,��2������Z�V�O˖�X��si�C>�dv�4��������	�}1��1�Tݫ���f ���UZ���/�a|�RN!�Q˜�\{�%�������=-�EEW��o��ú�Jx�}��h�%0зR~(�dɃO9��D��S�ym`�ф�y�W�TQ���9~Hs=,�yq��3TR����6>ĆB3]�@3�O3��L�e'�u�S����@�W����<: X�%�{_��G��_�Z������-f�45��'�"��sc;��4L$y#�uv"Zoڬ��g^zGب[:��E[ʍ�}��G,Z$r8�w"����0avbYn1��=�r,�L<�J �����:�sO��?�S�%H����~�||�KXM}�*"z��#���7֒\�M֠�]ɃE?y׈'���|���$;��IH�bj�10��s�t�zxsS���n ����e�"S
c�aV�g�I��)_̚%��Դ�U��xG&'�z�hg�D��In��W���R��1VO^��!{�7�,-��?�װ#���^�+	��߄6����3���^������:ڿ�gX���z�<4�ָ����όTl;�A����r=�͟���"�#D��j�?�����"E�ȡ�I���/�T?K�=�R�*Va�4�bHx��I���9��C���<��iiE`w<<\�m�'a?+��Z��y�v����~Rf�C9Z�r<p<�E4?&���p)f����8}��p��ބE.᭔��]�#�/�zs𐝨<��,����D>��Մ�.�Qq�݊|����(�E���
�$z2�?/��0P��wt��;��ջB��5	�Þ/�5�{J�������P��d2e#�lG8��"��@)�o+�&h���ߡ*q�|de]�V�D���3MS���F�����P^�M�Ϟ���q뮚�3R����N|9Jɂz�pB�s��u��4=�C���F?y8;:(_�'9W<h.��ih�8�RRXM��kZ��<3��\*��bmN�\�ϷG >w\���<���~X�·E07٤���[*6�O��q�Ѫ���=�`LD���	ߺV9�:�)%�`!���bV����"�8�^z��"<~����]@��)��o�$������_D ��qq&>�S��o�YG��W��t�|�!϶$4�"�lW�v�E��R���Y7�:Ҟ�U��S�
�!���(&�������Ӧ�ņ�A�8Ы�#�$�Sǁ.l\�|�� �lܗ�f(�"8�x#t��[��_����!q��Pw�l �п�H �Հ����Cv�
��[癃����N�>��4�i��_90%�f��V�g�lݓ�S)�p��:KQՉ"/��/8 @^_�ww���G��?�IsJ���
dQ��4�>����㙜�Wu�(���U�-HJ��"��S����EM��B�';H�� �#��3�#Zpi����ս�F|P�19D����_�_׏Z:냻��=��"u�}�cIiDH�4Q���A����h���tYF��u���6�8��4���#��Hu鵾�/x&Z|vf��Y-|�G���P�Zm�Xq�(�>�2B�N8�����Ls��o�"!�Tʨ����T�~��D��b!��b�X<��*������K/��n�@�>��+3U�q���?��FdiR�75����EҊ�l���oa�w�4łk�Y=��#�����zj�Ţ��+̭�gl�R�t��J��W(v���8.É�C �M��k��T1�W��``-�'�#&-"�!�x��X����JO�������\���P�w7[8@�� ��[���ƨѫh`X���ܸʦ9u?0�2R��O%nQ���֮�9c�Jx�te��.�ັ$ώ�/����-˦~+U�@XL�(��Ƿ@�d�/ ����l���Tq����4�:��E�w���⭇G�*�C�|�ȾM�(����Z�)��}�.=T	�&	P׻o7�v����M�f���5I�g�)�U3G^Ð-���v�������Y���@KF���k;*����ؚͿ��SH�����t���bT,,��>E�0�P?b�X+-b�Id��"K,�b�4s�_x�Q�����PK�r�N��WCfi����Nc~y�n7o�0��'��!|���*_t�Z5���_N��Ix)=<kK�czH	�����u����n�vW-�۸٫�jr����z�	�I%�>�K���<���b��9�+��镨��_��v|��	�\m3l�>-���8��IY������?�9ů�%Z��#�~Ż&ͻ�q6Y�:²k�b����u��E�S�64$C����>�!�uro~�XWI����!1r�݄� �i�é>?�Y�<z
�3+��_3��d��.uUס���8����{k���n�qZ��!��Pg�|��?��/��	�	���nn��"X�h<�q�`������D�Α"N�`�qzj&��J���t�1��`^.~,�ܔ�t�>��_75׏ ����{� 6O>z���fUv�.ϏS����ӏשs�Y<R5�+WMy i{��ݴp�e��y���]�!J�9::�		�̫!��0�cG-7��;�J_��u~}ݩ[�\xi��~T7�-�D,?�Lh�������ڙYC�:a%�ll�c��s�:
�-�������vЮT�F����� ��x��䐺$j^��.����]R@�-�N��\)�e�/t�m��˝x��\v�B��7ׂZ��=!$��4p���Oގl�Ţ`oD)��ˍ��GU^�Y�H��~���=:��su2��k���p�8��S?,�8�Z�H��	��	���2���#W^إ���ZA���D�" .T���34�e���������ӛǟ���K��,���m�M��e9I��i�Y��^~F��ԫ�ȹ%'��c�(W����+�<�E k�I�g���.��Gք���~y]�����ZD�Q�:�NH����oyţ�ುN�o���{[W5X8j�``v�]gk�ɣ�vͿ���ח9�ۙ[)V��l�xB��5Q$��tA+pX$G���S_����f{�n��i�zyjL�yPS�ݥ�z��@�ܢ&w��#�*t�\�@&��\`t$�_vx\ �(�p��aUu��x�}}{ݚ�����e�&��[�p6����0��5���LM�j�8��AR��`�$�9�ˡ.��ax f����t�h�c�>���9;\���q�����R��d����bk�����ⴧ���%�Z�98��4����\Di��1(s2��B�Q�6C�"�N�*�����O��m���X���z��Q4"���,��N��=���g/���9{���b�;8&ԁ0�Z2'54;ѡ���h��E8)~<'���s�_G���g����4$%p��H���'��-����uV�̴�H>��	�)�)��u�X��LйO�#^��-bߎ���[VD�#��q(�7V:5��C�J5������zF>�H��C���]/s��d��-(�~��u��#!4�.�@�v��8�7�97��G44I ���'ЊZ��2����]Q1�^5X+�c�N���zk�����廍����%~8	;�!rai�аhR�.����ǐ��v��;tp�����������=�=p���@�w�l�<�#��C��u����F:�e|����;
so�?=��Pֱ�]dl��������o�Eο-C�*�921�	P��l��EQ�]仐i�W���\��Ҧ���D�1�Ԅ<��Wֳ�ێ..f�@_w�E��Z��r��jP-����G�(�H*P�)�\���<�123�����t��u�:�\��2�����0y�^j��E$E��<UܽTEx@^�/f]u/��ّ��.�ޒB$���/kG��΁�x�q^ћ����h@��3�鲌�(���򉤒��
,�<�a�
���G�����O��Ȯ�k'N�4�03�L3��S����xa6L�<B�h��9q�5�u-�fI��S�_��$��Q�'�d���N�X>#���za�Rv��LF5v�)��:��)�Կ��sD���
ݥ6�~hL/���K�M}�lي)�����-��G���5M�䐉*]>����D�3aV�:UT �,��퇖���֓^��Ƹ�8  �>RvD�q��H�Swxo�,�^�K�8�&�	��xid����.���,y�����feZ�� h�YC:~/�c��
$�b���;C���
���-�"2����Ijt�K�5WF�!��>��qV�W*�Χ��J����,6u���!B%K�1������7�s�^}Ժ᰸wv�P��O���ر3�HR2$�7i��	��> �-~�o^�*b��ECPO���(��x����ӟ?7{	\�d#>�{)�.!E9��t�:�5 ���j�l��}�*o�G�]s"����@I�f&�DR�:l��%�0�3�β�P;�M/��s���R�c�_���4��O�y����3��J`>���aa� ��xnYv�T��%-�^u6�[ko:1(9����f����H��ik����!r�g��VbNIF&0�B������_�یk���癣Bx'8C��>d�'���{��N��^���F��8ݳ��4��E���t[-�Kc]5��]X��x��q6l�[%߹DCpV*�UU���%F�
A��ǅ��'��~��0L�4������j=B��L2������Y�͡
]2������-�L8��_SNƮ�!�y�p5R"r�1S�p�O��CM�������RϿ"���m���F0贒�g�5@��0��X����l=>`�hRLE=ri��8e�
Ǖؕ�oy�O�L ,�_��!7<.�'%���ޱ6w�=����3b��;��ε��o��~�=�C��M��z��3��A�:���h�l��^����XVuf8�S�CQ)6�N�Co���$��� ���Z�����U銛CH= ���W�RRR8a 1�5�q�gG3�$	�=>e@�
�Z� �`K�7��Wأ��pa��xnv��d���<�����t�Zg���W9�ޤ���`�jK�ں��X�@���+�kz�>����{��A��њdz����ٵ
�ܿOr}u~�:�T�w�&�51/[jBȲ�N���l��g7������W���&S��hv���߿GT_�~}4o�̉��_�� 3�\ҋ�e����{���"��$rY��?ŽX#O������yH�~6S���{������"cN]�!�ܦ����6 xXU3Z�g�H�5���1 ����
�l����i&����%5n�uKiADezm�J#���U������7�U@h��7'���$���D����������{�ŎǦ!f�H�#ֆ'm��+���Ki����r.��S�F�3�g��'���Q�|�k��M�K�a�Ey�����a���sp��{�f����L�T���
9P8~BM��	����i�L70q1�c���G��K������'+��#���<���4��݂1q�����wc��/7���b�B7�1PAjyj�C��-a&���P�j�\��]V__L�x#��4��+���/M����g�ZS�F����hM�x�J�9˧H��x�b3*��j&X��]�yH��,2V���W��:%F>�c�c̎��ؼe��!.hCմ�E��v�x���;a4Rh�+NY�#u����>CzۓZ��Âa]��=�q�˪�������j��N(��U��灖�N���F`UIՔ�u�Q�&N�#��'��S<��H.���dJ��3�XX��-��ۆ�a�|��{U����>^�N����D�������/�ڊ3Lޭ&^��Nyׇ�3�'���BR� pɇ�le����ܿ(�3=���6e@��;U�xemr�C�˟�M<$xw*�ی0�@��K�(�<;���ݕ�Z�f��-�q���S��6TT�GϹ@��r����\a�{Q��Z����?�J��ێo�~}�A��*+6���߄;3��B>R�P��o�9Ei��ɁvU�9dV��
�O�Ѐ����UxY ��T3e��m����t��t�Οj���E2r;r���k��&�+R�<D�ʼ==�����t���c�����e=Q�z��}\
�}�=BI��n/�>l?��f���c��5�xSo�.k����~�,B_G���R�����jn���wۜl��tu�Q�VуUJHL���FW�e�$�)KM#���%����� �������L�YG��H�\֬�D�k�>`�}�4R����Ǳ�'�#f(��cTş6�|}�U�يݨ�X@�VZY\�鋆� �LQm=�tk��O_��CO��u�-q�Fߎm�X�I��O1�ȬJ��ն��O2i��r��5��W�^lc#��O�	�P���.�7�z��C�f���L��O,R�4+g+S${6��!�;ht�y%ɿ���*+�@��J��5����f0@?ly��*�1^���gք8�m���,}�bҠω�%��T��:�3a)y����S�/��?#�� ��`
k�L��A������tgSǎd��@��#y����)���4�و���沁�=���'FE*վB��GzF�c��B%U�ơ{��pRN�S����)��=y�5�Bl��M��n�*�aS�h4��o�����·/*+f� ��0�~e=��*��,�(u��i�H����v���+���F�h��+^��^�f�@�y�g��>�{�Ր�IUE�����<��ll�,\P~	���|��|p�ɒ�bN�d��l��lj=�,"�rʥSm7�z �l�2�ɭ�z\�.`b-{$\S5�j�2iн��	���N�OR���K�o��P[����*��]aٯd׬��=-���D�c��t�W�?I4B>���Z�`t��w6}\��9�[� 5��P*�����.��8 ���2��iJ���
���2�����'��X��>'��� XB&A��X���)Z�B������T,��m�&�j�ֽُ�Q���4���AKw�%/|l����S7��0k���[�W������w�GQ����ܥ�U���&b6�7d���5}�����$�/��K��9μ�G�.ϯ�9^�z¾�Uy_����y����f|MOb�Y�̲�$O��Ŗ܃�w�M5�5��1m����~��k>%�b �pA2 �?�I���� �$�j�74tYE�K�LA[@\&Ԗm�B!;�7/q��
uǇ���I����h�f�';� Fb�6ֹ},(�K��o���G���Nv��%\<mq�<��E�t1k��P��R��BQ/�*��z���		�P����"�$>��Բ��i�*ly�ђ;e&�ER��B�%���¿�o�N�zC1��E�z�� �'`)�<vx}[B34:)��7�b"
�!��R�9'7D��l��e�����'�(h���%�ǂvc3R`V��BW��zª1�-#���зX^Y^��U����q�S��9��s�6����������@�X����-�^�]Ґ:/Dddʌ3��.�=�J�f}|�{�>M���=4��	���jT�ŷ�x�, �J^aA �Ӏ%�HNn�E�~���~���x|�r�Y��3�����-�d��.:����Y�QIx��ep�VI!`@�![�x��b��\��$��A�[�/� M�GȬ[�|p>���73�u��e����y�W3������}�������n2���V%fw�\�A��#[yXI�&C���c��I]�~p��?C��t�'MKY�m�t�:*����tL%�A��<��J���ݕâuًdxQ%�莇��:]}����J����X	�5_�����.Z<Hd^���%8G1�cl�,��5
��т
U�#�c�W���r��h>u������n>y�F��AU�n���$�I��i/f��Y�D�����0��@u`EDg��f)&��p[ ��F�5��h�Wgx��>�1�<�J����3C�z�-��"��O�R<�RR�Ӟ:��p�>�):��L��7�)����]�w��p�:�Я.��i�r_�+#jWN�}ӥA'�l�l�ex�oYH��խW7���3�<��r!������R���P�{s·�HI�tzT2�uM�$�\�-l7ر�N�H[X�KJ r;��xnb{�UFv�XYY��Z������%Xp[��Q4B���a�нI����$2`<*�B>|���W��!���i)C�ZZ�~M��h��u,(S6*Q@l��f�e��P��R3�#"�������� �-"�+�/�v^���sj*��j	��q]�������~�s��2��"�!�;װ�E����	aF�*�#�o��o�`~��� Z�H��J)*w28������y\��֚B�2�x��Yj{%Km-�]�T��5vg�1��q�4!.���8!�!���E4&�� 8s0�~�Z�UN�ç1�{�rM���TkXks�"H8<$�W�� �=?����S�Y����:����q^�t'��%�'��u�� �l��@��a�sֿ~�T >IR�����<��!m��?XU��E�q�`�A��RtV�P�s��;���;�;�I�s��� ������x����R�BfF���rNf!Q2���c:Fه��*�콎Q�ٛ�s�u�8�������s����w�����|��u]�+�hЙ�2������c�ᗍ��aʨA_�T��;�v� PF��9�OU�=Ëv"/�9�'�)_`��Ű��ޮ��c�rw�w�mu�+�
��X��g9a�Z��ݷ�oB�TG��������2vʦG���ۻϡ7+&Z�y	�5��=�9	��
��nm�)�LΛ� ���M�ؾWl���Y�s�
zc���'���d�M&�Z6��NfX��Eċm"�����S�Z�hF���mV(��	�JN�{�p���R� ��~x��"eEcqqq�H�4���1�ҝyKq�OO��N�������֝�t�ҁ�lT�X�1j����)���s��$PL)���@X� ���	ٸhמ]'d�B�/(�*`�N�*��_��};���d�Y)¡Ĝ��Pt�ɔ�3����Ao�T���d�8N�h�ED��ᗛ�'%������T�M>�{��*��H{7�wF,���q�����������?�ѠM5�_Bӱy�5�&��_`8$�o�`�J�<:-��f�$��b�� �?����xle�)���â�0!�_ƨ��)|r�W�m������Q��^;Mb{�To���)d3[v�U�W8�i�b�sEχh@���׼� 0����U]-�C��Ĵ]6�Y�����|fgsMP� ��L���ݾ�>�,�M5�n�56�.-}5M� ���,,���r
�N[_�e�or����U
����&�,�-���A{�y�jA`Ư��/���`�*�a6b�T;'w���&�/�R��*�M/�4��:���\M3��1?�-��T���XV�v$���Af��>Rl�e�w�W(⼁�K��������X�;'������&� {9�S��upk̴e~��B��o3-Ѵ4�?%��o��Qj3�]<ɱ���%�~�^r����2����lo	�m�f�Wnw��J;p+3��&Q�_q�����@�n��e
�ZqZ�]/;PȜ~�r��~	)��tշ l����C���|vx
���u̫�&����K�y�࿳%,�$���t����5'�f[��|����37����Fw�'ؠo���*�Lt:���m��=����[0%�]WU-!�%�����Cń�EyDy�<fpX������lϜ����%���p��6�	�຺VR����ln�`���S�#�j����k���y�2y^�w���ҝD�\A���Ďy�u�q�w��WD��5��@��2���n5+^��l0����=P7��i���Z����uE�T�o`	s��}��@��F�H��2k�BO3��k�Sʢ��u�YB�Xg��rd� (��{��:������,U'R�R��C��Y+n�ǥ�	Fn����e�3Y,��,��˦r.Į%V`�z$�=yh�)A�hɽi��߈i	��F�^���dд�'��Bt��{���$[���f�g�b�hk��ߏ��~�a
������Fk��r�8�;F�T@0w�j.�T����C�1���WrYl�܊��Dx��%�=<�Т��l�+^�e�XwY�/�ȥ��S`� ���g6�����w�E����ߤ�޾	b�a�v��`��ǜ���>�@��ojS�L@�"��LPX������8�����|��ٯ1�θB���tC�s��N"敉B;��qY����p��<��t����rJD��fL%��&b���0/P#�\��>������_Ks�+�v7�oz�,�׼Eʩp�!�ﻤ��Y��ެ��-+h�<�9�gS�g�2�p�Gb.@=�X�-`>�j��Tc�����)���$sp�N��jZ�cRn (ۼv���=���X5�^�x��I5�G
�0,����˹Sj��V`��]���Sƭ�>-�}|f�Zl�j��_ѳ��e�i�>y�G��/A?�ػ�����f�	c'��τY@-��7�,�43Eⴷ�R�,oH��M�ʹ��0�xܾm1S��Fy'�B9��W;}���^����{�Ɖ)-"�L=x1�=gS�<����/��T']BƵA���"Y&hݴħ�?��T�
��rE^��.�̸�nۑV�,/��Я�W�(ߠ��u������R�.�ݺySGp�Y4�U[�$	��Y��
�:�7P0� i2+���+s,p;Mt�!J4���LxMܯ@��/R��%��Í�RG��YTU^UV���&��q��>Ck~~	����T#��(����c�ۉ~͆��T�����C�^��%.�&�b��<��B�*ޢ�r�rxTd��iz��VB���\_�u���N^��{�_�Z�2`��w[N�M��o5)p�Mۘ	��o����GD��gϑ�/��c����Ί��K���tj��O��S$bo���N;D��z�W�ơ�?�I�8ؚr��)-]��%�Vt�j���Q�����i��p������o��@���j�jD�|�s\���z0�fQӁ�D��D���0;4�Cҏ�=ن�A���p�O�QD����{���.NS!Q�� ƓL8���GqQi����6��
ucs3�������E�DA�LW�$*�%j��/���~t��wTkN�L��:5��P��iUPo���R��=�4q��\I`ҵ�7��f��� �b�>���㲴��48x5o��0�#K����g�cE0f&�wr�\nQ��>�_������r�����Y͗90���y�3����I��t,j^-�uZ �0,��)c�D���B�8y�\�8�K��p����+*��q�JoQQ��Ѝd�р8v���f�=흋��0�zM	A7m��|����<�UO!����^�J4��q#�>�������_k��n���];P����z�X�����!�=�stړ���š:7�����|�Pg��):8�r��S��=��9��Ҷ��iJ��P:0�����Ga)Li����u0���'{ZZ�����9���.�
�25JB���
��ӆ�>��i�V�R���G��^���!�^�NW�k^nw:�?�3���iCkK��K<eC�h*n��6in5r��p_�EC��Sx��+w�ءkC�4�N�
��ŕ�:R��i@]��Cu���,K4���7��\�dM=n�c:}���%c������<�@`A�Y�gZ���].�"�ˏ��k
'e	`諣�]"^�?�ϱ��l��� cPK��l����)�Dno[ZZ2 ������C������d�l����5P�k!�I�<��y�\}��?�X��T��13�m�������y�� +L�nM�_��M����@Rv�d�FP�r��;r�+g��á��=[c*��z�����+��@2���*՞�I_[�;�qR���ցtIb�(�N�%��8T��_�I����<C�����XD�����ȼŞ�
�짻������.	��p����4�����Ki���N3-�x�m���g��d��P	��d�h4UѨb��bhg�����ү<Z�Uq�Qs�ڟ����^710�9����\�6[�y���5��v��ٱ��Ɉ�����T;��hQ��Y���#T4�>e�ҊC_���{�%�rϯ�
�$'qk��Q�$=vs��[�]��N��p�n�Y<z>��i�`���jZ'�кA��)�D�y%���qL������`�q2�G��<���׋��Rs��<��>�G:�Խr`h�B�D"z���)��Z {�����L*G�
��������#��ff�����р��Zq'���K�[�EM�Ϯ��3&�,ƣ?]�<w�O0�S�?��o��F�l���|A��� �%<d�ݜ�jJ>�R;�-�A���x�'��� @�׆�,�E�ڄ+dt}���}��"�mo�&$D;�[��.i^�)�q�D��`'�A8��m�{ytڷa�ɝ��̘�V��-ZDNB�mDW_3K��M��V� �x~O��xHȟ��s6EҢ޷�W��R�W��� �|`	ʮ����t*0�ֻ����ơ[��r����ZH�O�4�%;g#�ڱ
8>+;MK[F�w���Ap�#�5��Z�&��n�x�~���M�pʺ���tg����}�s��׷��>۝��h����mM�TD,֘l�y����t��ԴW���ڵљ�j3���zd{w�B�u�h uoDr�9P.D�ã��j��H�w��hm?q�[������d�6�<Z��o�C�摮Hl ��S�OW�{1�#�0���̅�1Ou	~�L���ή�[��c�G{Y��C��GG�|ȶ)��?_�u9SW�1���/i_�q$%��n������	�ɗ��7s2[{����j�K�<�4��iC�DV`<�\	�
!�G�wb�\'%u�h~�:.ì�����`].m��He��i(L��T�>�N�,��V/Oh�:�B�E�bv��m�o�m��>�y�$��v���f��xooo@
0K�A�4��L���Ņ8Fʷ}Fky�K�E�K<���N]ԁ���`�D���E�k��~~�l���T&���L�U�ޫ5�H��y��o���^���v��V����f~���z'�V,�p�`�19oA:�۸��x��I[�K=�{%�{�tv^m���U܎eI���w~�xSSSM@�5E����O��V��[)��O0(,��ni�:��,W,&���f[��)������Ύ��4�q�Ä��Y��_����z��<�	�5Rm�L����)�_���	̲D��ؼ���77��ģxOZJ��<�,��~^Ps�FV�;/vCS~ƣ�k�_q�؝����7�-υ,�8h��x����ư((��PK8r.�=�ݝ�x�>+x�z�jh�z�b�{i����oMU5ǰ�DL���Nfk�A
zJ1>Vؤ�i��S8�D�c��#�7�L*����U��8a�7'�KH°8�?<M�x���� �iD(���W�<V]�_%|�	q�g�ޣ́���{�˄���.�h'�T��r�w�����;�������.6��v��=�F�=n%+Ϗ^9i����B���l�zrr+�x_�}A�m6���վCvbvvz���"Hi�A���r �'?5x_H���I�B;���`�}��Z��H򷛖槐���u��b�u�r��4�7��Ji�5��� �̕�cξ����]��ZA��mki��>���x���Y���S�2��q�	���2�v&K�����k���i���4g��^�k��?%V��@�`�,���q&i}��=q�`�� �_��K��%"���}I�,O�x�8K��tM(!���+qMMM����wzFdqA�?��zO��3,�}��˦ކ�@���Q^?�5�Ot��]����2N��\p�|R]�KeSWt���[B���z��������G�+�����2��N�P<1�̗.>9�.ra�[ꪜ_*w��&#ݛ�U%�V�7�e��-;��������o���w6�K�njUPOkh�3<{n|��r��ur0;�����a�;G�׵zŖN���!�ٿd�N��R���[�����JJ&+<�`���.��-߆�����>����.��ZU� =O��Է�,v`=���wrZ���%^��xuϰ��רHl �0��_^}��K�d�J�\�Bԯ�.[�0є�0_B���m�R�õ9I�s��M5s}F�p�3�����}��q�m��IU�n�p��yBxr'���LL��ۼ�@�y"��K+=�����Yi.��u����7�p���_Ml H����}��)ݟ�W�R��\�ܧ��}��+�a��u%��݅4ю��^7��e��h\VK\{,�/٭#V�gw�Tm�m����YQ��}�
� �70`>�p�o��%�O�E�\�+��jBR���#OUth����!��lwǡ����-] ��
�
Cx�#5f�_����)�0�������'S�������G׽bW��(�hs"�ד�&=-�1k��W����'(,�ə0N�~(b����\h9+��\3�3Z��$
*(�\�[��q��%t۶�q�.�^�q��F8�Ou{G�$:�W~�X�.X�G�rf����8�o�A��{#zgb�ls�ޝ�Q?�8���[���1c�#�=čO]�+��:-n���VY\��[�о�3��մ��ƞ�������T,M֊&�������c�k��ג���T��˄��Y(c�UC�dBc1�p��.I�<��fȗhW2��_G9*-�}�"B�Kd�E�l ��搏
���n�SI7�h���(Y�d���o�9g\�j��`¸9��Էr&*�)2�M�7��}?! R����8�;_�����[��d�l�f�,Γ �G�K����h�Ϗ�#�M1�*��J0v2�ˢ^����&���s��k�{җ�ֹ�ls�|K{ѫ%����� ��5	�(ƀm!�#+>'�TG�Ѕo�a�L{���x���k��1������eo��s{�A�ʒd�%4*�1��� �ޟ�/۴vVt��Q=K�hj�B�1�s-A�/^E'��Y�ٚ�?�X����lyC�.sH������t�v����(���3��&�񇞥�ty�Ct�� ��?�s5L|�k�4oGY�O��sp4��w|R��b~�q<����m�DP�|I{�R(����s����*pބ�v�;��i��n�`���J�&$A��9m��`���g��E�;�
 �#d(����`���n�'�WUa�?��7X�/�d���,����}�{����D��Aq���R�:R�Ó�6�5���!^S>W玵~h����а�L�����e��[��/Ѻm)�Q�s7�����x�x�`���C;|j[������ Y�x�S��@������+!�	c�V����9�y�썌j=l%���k���LR�(ü�hَ�\C�aok�z?֥,cm+z����t�1�Z�r��~��R@���*��Գ�=���v�A��w��J6����lR!���D��4&$��}p�����=ٳ�(��~"�� �:�c_�C�@��	�]R����0��̚�Q�1��.���vf�����#��U���t�kZ�g^~���8 ��2ļ�W�1��� �������@�b�?�"�2�x�R�ct��5�X�l���M
v��!m�gc�;�����"�,����R������~�+8ǣ�<�S���V�G;U�j�-����}��=Ԗ"�X�8�o��ø�U}B� :�řJ	�\�x��!D�F*��`~���0zb� �����1�ycF�u_�	30���#�VW�k�\�ABz:Nu�
7� �G�����x�%
�N��T$�k�2÷���TY��3v/�d�ž׌����|�Y����� ��`����@ǽf���~`����f�j�|��s�[�,Y(�gvq��q�9�K��k�� -BI��5}�b�%���0$u SYL�r�n�;�ʆW��J�p���i��ia�`pʙd���[��^s���}��� ȳ���5��Ҍ�Ţgfzk�Xk�P����?{ 	�y�P�w� P8�Ȭĸv��7 Dqi`sE��d#ms�s��Խ�Ѕ^�����{AL떑V�0�$�i_����}��?�������Ԥ�ҿR�<W<�L� ̯9y�ބB�~<w{;����E
tG��6�G<��xTv�%�a��t�2�R�~�4&���/	>��;�X�;��N��g{��J:�v�>!��|3�>�6j!P����DT ]2^�7�e�/�Y���_��X.�����?�¸|xi�C��?�?PK   G�~S��ME�  �     jsons/user_defined.json�Ok�0ſJ�96�%�OnKs	tKi��%��G�JvK��%MMa�]z������捴%��2%C �@�L��`��Mi��IV�5������Z�����ʋţ�6J�Ã�l$��z1{�.'ĨHT e"��S.�ZiH�:�$�L�DNtt�N{?����ƛ�?<y�1�H|���u�έvd�%vX�L�Z��t-Ir�
����S��=�k4e���#Y��Y>��wx�]�7��bg?ir7y����X�ΏI���F���*�Z�֙Lʬ�r�u�s�i���H��)�^��rL�������Ђ��E��1�����N�6��i�X�'eY�U��=&��ͣ�>���D�>�������%nj<?����
�����~�_����PK
   G�~S�8��  �.                  cirkitFile.jsonPK
   ؚ~Sk2��XP  �Q  /             �  images/0deaa9e5-55e1-404a-9dfe-2921a303d637.pngPK
   g�~S��RC�c  q  /             hm  images/e1605cfb-dd4b-4fdf-9f1a-7191204fc245.pngPK
   G�~S��ME�  �               <�  jsons/user_defined.jsonPK      <  ��    